`define NFLOOR 10 //Number of floors in the building